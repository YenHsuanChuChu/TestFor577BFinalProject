`timescale 1ns/10ps
`include "./design/Pipeline.v"

module cmp16 (
    input clk, input reset,
    input [0:31]node0_inst_in,
    input [0:63]node0_d_in,
    output [0:31] node0_pc_out,
    output [0:63] node0_d_out,
    output [0:31] node0_addr_out,
    output node0_memWrEn,
    output node0_memEn,
    output [0:1] node0_addr_nic,
    output [0:63] node0_din_nic,
    input [0:63] node0_dout_nic,
    output node0_nicEn,
    output node0_nicWrEn,

    input [0:31]node1_inst_in,
    input [0:63]node1_d_in,
    output [0:31] node1_pc_out,
    output [0:63] node1_d_out,
    output [0:31] node1_addr_out,
    output node1_memWrEn,
    output node1_memEn,
    output [0:1] node1_addr_nic,
    output [0:63] node1_din_nic,
    input [0:63] node1_dout_nic,
    output node1_nicEn,
    output node1_nicWrEn,

    input [0:31]node2_inst_in,
    input [0:63]node2_d_in,
    output [0:31] node2_pc_out,
    output [0:63] node2_d_out,
    output [0:31] node2_addr_out,
    output node2_memWrEn,
    output node2_memEn,
    output [0:1] node2_addr_nic,
    output [0:63] node2_din_nic,
    input [0:63] node2_dout_nic,
    output node2_nicEn,
    output node2_nicWrEn,

    input [0:31]node3_inst_in,
    input [0:63]node3_d_in,
    output [0:31] node3_pc_out,
    output [0:63] node3_d_out,
    output [0:31] node3_addr_out,
    output node3_memWrEn,
    output node3_memEn,
    output [0:1] node3_addr_nic,
    output [0:63] node3_din_nic,
    input [0:63] node3_dout_nic,
    output node3_nicEn,
    output node3_nicWrEn,

    input [0:31]node4_inst_in,
    input [0:63]node4_d_in,
    output [0:31] node4_pc_out,
    output [0:63] node4_d_out,
    output [0:31] node4_addr_out,
    output node4_memWrEn,
    output node4_memEn,
    output [0:1] node4_addr_nic,
    output [0:63] node4_din_nic,
    input [0:63] node4_dout_nic,
    output node4_nicEn,
    output node4_nicWrEn,

    input [0:31]node5_inst_in,
    input [0:63]node5_d_in,
    output [0:31] node5_pc_out,
    output [0:63] node5_d_out,
    output [0:31] node5_addr_out,
    output node5_memWrEn,
    output node5_memEn,
    output [0:1] node5_addr_nic,
    output [0:63] node5_din_nic,
    input [0:63] node5_dout_nic,
    output node5_nicEn,
    output node5_nicWrEn,

    input [0:31]node6_inst_in,
    input [0:63]node6_d_in,
    output [0:31] node6_pc_out,
    output [0:63] node6_d_out,
    output [0:31] node6_addr_out,
    output node6_memWrEn,
    output node6_memEn,
    output [0:1] node6_addr_nic,
    output [0:63] node6_din_nic,
    input [0:63] node6_dout_nic,
    output node6_nicEn,
    output node6_nicWrEn,

    input [0:31]node7_inst_in,
    input [0:63]node7_d_in,
    output [0:31] node7_pc_out,
    output [0:63] node7_d_out,
    output [0:31] node7_addr_out,
    output node7_memWrEn,
    output node7_memEn,
    output [0:1] node7_addr_nic,
    output [0:63] node7_din_nic,
    input [0:63] node7_dout_nic,
    output node7_nicEn,
    output node7_nicWrEn,

    input [0:31]node8_inst_in,
    input [0:63]node8_d_in,
    output [0:31] node8_pc_out,
    output [0:63] node8_d_out,
    output [0:31] node8_addr_out,
    output node8_memWrEn,
    output node8_memEn,
    output [0:1] node8_addr_nic,
    output [0:63] node8_din_nic,
    input [0:63] node8_dout_nic,
    output node8_nicEn,
    output node8_nicWrEn,

    input [0:31]node9_inst_in,
    input [0:63]node9_d_in,
    output [0:31] node9_pc_out,
    output [0:63] node9_d_out,
    output [0:31] node9_addr_out,
    output node9_memWrEn,
    output node9_memEn,
    output [0:1] node9_addr_nic,
    output [0:63] node9_din_nic,
    input [0:63] node9_dout_nic,
    output node9_nicEn,
    output node9_nicWrEn,

    input [0:31]node10_inst_in,
    input [0:63]node10_d_in,
    output [0:31] node10_pc_out,
    output [0:63] node10_d_out,
    output [0:31] node10_addr_out,
    output node10_memWrEn,
    output node10_memEn,
    output [0:1] node10_addr_nic,
    output [0:63] node10_din_nic,
    input [0:63] node10_dout_nic,
    output node10_nicEn,
    output node10_nicWrEn,

    input [0:31]node11_inst_in,
    input [0:63]node11_d_in,
    output [0:31] node11_pc_out,
    output [0:63] node11_d_out,
    output [0:31] node11_addr_out,
    output node11_memWrEn,
    output node11_memEn,
    output [0:1] node11_addr_nic,
    output [0:63] node11_din_nic,
    input [0:63] node11_dout_nic,
    output node11_nicEn,
    output node11_nicWrEn,

    input [0:31]node12_inst_in,
    input [0:63]node12_d_in,
    output [0:31] node12_pc_out,
    output [0:63] node12_d_out,
    output [0:31] node12_addr_out,
    output node12_memWrEn,
    output node12_memEn,
    output [0:1] node12_addr_nic,
    output [0:63] node12_din_nic,
    input [0:63] node12_dout_nic,
    output node12_nicEn,
    output node12_nicWrEn,

    input [0:31]node13_inst_in,
    input [0:63]node13_d_in,
    output [0:31] node13_pc_out,
    output [0:63] node13_d_out,
    output [0:31] node13_addr_out,
    output node13_memWrEn,
    output node13_memEn,
    output [0:1] node13_addr_nic,
    output [0:63] node13_din_nic,
    input [0:63] node13_dout_nic,
    output node13_nicEn,
    output node13_nicWrEn,

    input [0:31]node14_inst_in,
    input [0:63]node14_d_in,
    output [0:31] node14_pc_out,
    output [0:63] node14_d_out,
    output [0:31] node14_addr_out,
    output node14_memWrEn,
    output node14_memEn,
    output [0:1] node14_addr_nic,
    output [0:63] node14_din_nic,
    input [0:63] node14_dout_nic,
    output node14_nicEn,
    output node14_nicWrEn,

    input [0:31]node15_inst_in,
    input [0:63]node15_d_in,
    output [0:31] node15_pc_out,
    output [0:63] node15_d_out,
    output [0:31] node15_addr_out,
    output node15_memWrEn,
    output node15_memEn,
    output [0:1] node15_addr_nic,
    output [0:63] node15_din_nic,
    input [0:63] node15_dout_nic,
    output node15_nicEn,
    output node15_nicWrEn
);

  TOP pipeline_node0 (.clk(clk), .reset(reset), .Instr_from_imem(node0_inst_in), .PC(node0_pc_out), .memEn_to_dmem(node0_memEn), .memWrEn_to_dmem(node0_memWrEn), .memAddr_to_dmem(node0_addr_out), .data_to_dmem(node0_d_out), .data_from_dmem(node0_d_in), .addr_nic(node0_addr_nic), .din_to_nic(node0_din_nic), .dout_from_nic(node0_dout_nic), .nicEn(node0_nicEn), .nicWrEn(node0_nicWrEn));
  TOP pipeline_node1 (.clk(clk), .reset(reset), .Instr_from_imem(node1_inst_in), .PC(node1_pc_out), .memEn_to_dmem(node1_memEn), .memWrEn_to_dmem(node1_memWrEn), .memAddr_to_dmem(node1_addr_out), .data_to_dmem(node1_d_out), .data_from_dmem(node1_d_in), .addr_nic(node1_addr_nic), .din_to_nic(node1_din_nic), .dout_from_nic(node1_dout_nic), .nicEn(node1_nicEn), .nicWrEn(node1_nicWrEn));
  TOP pipeline_node2 (.clk(clk), .reset(reset), .Instr_from_imem(node2_inst_in), .PC(node2_pc_out), .memEn_to_dmem(node2_memEn), .memWrEn_to_dmem(node2_memWrEn), .memAddr_to_dmem(node2_addr_out), .data_to_dmem(node2_d_out), .data_from_dmem(node2_d_in), .addr_nic(node2_addr_nic), .din_to_nic(node2_din_nic), .dout_from_nic(node2_dout_nic), .nicEn(node2_nicEn), .nicWrEn(node2_nicWrEn));
  TOP pipeline_node3 (.clk(clk), .reset(reset), .Instr_from_imem(node3_inst_in), .PC(node3_pc_out), .memEn_to_dmem(node3_memEn), .memWrEn_to_dmem(node3_memWrEn), .memAddr_to_dmem(node3_addr_out), .data_to_dmem(node3_d_out), .data_from_dmem(node3_d_in), .addr_nic(node3_addr_nic), .din_to_nic(node3_din_nic), .dout_from_nic(node3_dout_nic), .nicEn(node3_nicEn), .nicWrEn(node3_nicWrEn));
  TOP pipeline_node4 (.clk(clk), .reset(reset), .Instr_from_imem(node4_inst_in), .PC(node4_pc_out), .memEn_to_dmem(node4_memEn), .memWrEn_to_dmem(node4_memWrEn), .memAddr_to_dmem(node4_addr_out), .data_to_dmem(node4_d_out), .data_from_dmem(node4_d_in), .addr_nic(node4_addr_nic), .din_to_nic(node4_din_nic), .dout_from_nic(node4_dout_nic), .nicEn(node4_nicEn), .nicWrEn(node4_nicWrEn));
  TOP pipeline_node5 (.clk(clk), .reset(reset), .Instr_from_imem(node5_inst_in), .PC(node5_pc_out), .memEn_to_dmem(node5_memEn), .memWrEn_to_dmem(node5_memWrEn), .memAddr_to_dmem(node5_addr_out), .data_to_dmem(node5_d_out), .data_from_dmem(node5_d_in), .addr_nic(node5_addr_nic), .din_to_nic(node5_din_nic), .dout_from_nic(node5_dout_nic), .nicEn(node5_nicEn), .nicWrEn(node5_nicWrEn));
  TOP pipeline_node6 (.clk(clk), .reset(reset), .Instr_from_imem(node6_inst_in), .PC(node6_pc_out), .memEn_to_dmem(node6_memEn), .memWrEn_to_dmem(node6_memWrEn), .memAddr_to_dmem(node6_addr_out), .data_to_dmem(node6_d_out), .data_from_dmem(node6_d_in), .addr_nic(node6_addr_nic), .din_to_nic(node6_din_nic), .dout_from_nic(node6_dout_nic), .nicEn(node6_nicEn), .nicWrEn(node6_nicWrEn));
  TOP pipeline_node7 (.clk(clk), .reset(reset), .Instr_from_imem(node7_inst_in), .PC(node7_pc_out), .memEn_to_dmem(node7_memEn), .memWrEn_to_dmem(node7_memWrEn), .memAddr_to_dmem(node7_addr_out), .data_to_dmem(node7_d_out), .data_from_dmem(node7_d_in), .addr_nic(node7_addr_nic), .din_to_nic(node7_din_nic), .dout_from_nic(node7_dout_nic), .nicEn(node7_nicEn), .nicWrEn(node7_nicWrEn));
  TOP pipeline_node8 (.clk(clk), .reset(reset), .Instr_from_imem(node8_inst_in), .PC(node8_pc_out), .memEn_to_dmem(node8_memEn), .memWrEn_to_dmem(node8_memWrEn), .memAddr_to_dmem(node8_addr_out), .data_to_dmem(node8_d_out), .data_from_dmem(node8_d_in), .addr_nic(node8_addr_nic), .din_to_nic(node8_din_nic), .dout_from_nic(node8_dout_nic), .nicEn(node8_nicEn), .nicWrEn(node8_nicWrEn));
  TOP pipeline_node9 (.clk(clk), .reset(reset), .Instr_from_imem(node9_inst_in), .PC(node9_pc_out), .memEn_to_dmem(node9_memEn), .memWrEn_to_dmem(node9_memWrEn), .memAddr_to_dmem(node9_addr_out), .data_to_dmem(node9_d_out), .data_from_dmem(node9_d_in), .addr_nic(node9_addr_nic), .din_to_nic(node9_din_nic), .dout_from_nic(node9_dout_nic), .nicEn(node9_nicEn), .nicWrEn(node9_nicWrEn));
  TOP pipeline_node10 (.clk(clk), .reset(reset), .Instr_from_imem(node10_inst_in), .PC(node10_pc_out), .memEn_to_dmem(node10_memEn), .memWrEn_to_dmem(node10_memWrEn), .memAddr_to_dmem(node10_addr_out), .data_to_dmem(node10_d_out), .data_from_dmem(node10_d_in), .addr_nic(node10_addr_nic), .din_to_nic(node10_din_nic), .dout_from_nic(node10_dout_nic), .nicEn(node10_nicEn), .nicWrEn(node10_nicWrEn));
  TOP pipeline_node11 (.clk(clk), .reset(reset), .Instr_from_imem(node11_inst_in), .PC(node11_pc_out), .memEn_to_dmem(node11_memEn), .memWrEn_to_dmem(node11_memWrEn), .memAddr_to_dmem(node11_addr_out), .data_to_dmem(node11_d_out), .data_from_dmem(node11_d_in), .addr_nic(node11_addr_nic), .din_to_nic(node11_din_nic), .dout_from_nic(node11_dout_nic), .nicEn(node11_nicEn), .nicWrEn(node11_nicWrEn));
  TOP pipeline_node12 (.clk(clk), .reset(reset), .Instr_from_imem(node12_inst_in), .PC(node12_pc_out), .memEn_to_dmem(node12_memEn), .memWrEn_to_dmem(node12_memWrEn), .memAddr_to_dmem(node12_addr_out), .data_to_dmem(node12_d_out), .data_from_dmem(node12_d_in), .addr_nic(node12_addr_nic), .din_to_nic(node12_din_nic), .dout_from_nic(node12_dout_nic), .nicEn(node12_nicEn), .nicWrEn(node12_nicWrEn));
  TOP pipeline_node13 (.clk(clk), .reset(reset), .Instr_from_imem(node13_inst_in), .PC(node13_pc_out), .memEn_to_dmem(node13_memEn), .memWrEn_to_dmem(node13_memWrEn), .memAddr_to_dmem(node13_addr_out), .data_to_dmem(node13_d_out), .data_from_dmem(node13_d_in), .addr_nic(node13_addr_nic), .din_to_nic(node13_din_nic), .dout_from_nic(node13_dout_nic), .nicEn(node13_nicEn), .nicWrEn(node13_nicWrEn));
  TOP pipeline_node14 (.clk(clk), .reset(reset), .Instr_from_imem(node14_inst_in), .PC(node14_pc_out), .memEn_to_dmem(node14_memEn), .memWrEn_to_dmem(node14_memWrEn), .memAddr_to_dmem(node14_addr_out), .data_to_dmem(node14_d_out), .data_from_dmem(node14_d_in), .addr_nic(node14_addr_nic), .din_to_nic(node14_din_nic), .dout_from_nic(node14_dout_nic), .nicEn(node14_nicEn), .nicWrEn(node14_nicWrEn));
  TOP pipeline_node15 (.clk(clk), .reset(reset), .Instr_from_imem(node15_inst_in), .PC(node15_pc_out), .memEn_to_dmem(node15_memEn), .memWrEn_to_dmem(node15_memWrEn), .memAddr_to_dmem(node15_addr_out), .data_to_dmem(node15_d_out), .data_from_dmem(node15_d_in), .addr_nic(node15_addr_nic), .din_to_nic(node15_din_nic), .dout_from_nic(node15_dout_nic), .nicEn(node15_nicEn), .nicWrEn(node15_nicWrEn));


endmodule



